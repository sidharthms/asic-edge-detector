// $Id: $
// File name:   ARM.sv
// Created:     4/26/2014
// Author:      Suppatach Sabpisal
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: ARM Processor

module ARM(
);
	//Nothing here
endmodule
