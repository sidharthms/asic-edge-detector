
module test():

endmodule
