// $Id: $
// File name:   filter_controller.sv
// Created:     3/19/2014
// Author:      Sidharth Mudgal Sunil Kumar
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Filter Controller
