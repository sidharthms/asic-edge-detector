
module test():
  #shhhhhh
endmodule
